.title KiCad schematic
C3 GND +3V3 22uF 10V
F1 Net-_D1-Pad1_ /VIN Fuse 24V/1A
C1 /VIN GND 0.1uF 50V
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ Diode 40V/3A
U2 GND +3V3 +5V 3.3V/1A
C2 +5V GND 22uF 10V
J1 Net-_D1-Pad2_ GND Power Input
U1 GND +5V /VIN 5V/1A
H2 M2_MountingHole
H3 M2_MountingHole
H4 M2_MountingHole
J2 +5V GND +3V3 GND /RO GND /DE_RE /DI Header 2x4P
R1 +5V Net-_D2-Pad2_ 220R
D2 GND Net-_D2-Pad2_ Blue LED
R8 /DI GND 10K
C5 +3V3 GND 10uF 10V
C4 +3V3 GND 0.1uF 50V
R3 /a1 +3V3 20K
J3 /b1 /a1 NC_01 /VDD /VDD NC_02 /VSS /VSS GND 8P8C
U3 /RO /DE_RE /DE_RE /DI GND /a1 /b1 +3V3 RS-485
R2 /RO +3V3 10K
R4 Net-_JP3-Pad1_ +3V3 4K7
JP3 Net-_JP3-Pad1_ /DE_RE drive EN
R6 /DE_RE GND 10K
JP1 GND /VSS GND EN
JP2 /VIN /VDD VIN EN
R7 /b1 GND 20K
R5 /a1 /b1 120R
TP2 GND TP_GND
TP1 /VIN TP_VIN
TP6 /DI TP_DI
TP7 /DE_RE TP_DE_RE
TP5 /RO TP_RO
TP4 +3V3 TP_3V3
TP3 +5V TP_5V
TP8 GND TP_GND
TP9 /a1 TP_A1
TP10 /b1 TP_B1
.end
